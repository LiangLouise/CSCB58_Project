

module Project_Banqi();

endmodule

module 



module initilize_game_board(ram);



endmodule


module control(clk, resetn, go);
	input clk, resetn, go;
	
	
	
endmodule


module datapath();
endmodule
